       "LR��\�Y�w���:����	]G��rIS[5   
<p>git klon git@github.com:user-tax/user.tax.git</p>    ϘÅ�i��c��#s�5�A'Sm�	y���n   <p>curl https://sh.rustup.rs -sSf | sh -s -- --default-verktygskedja varje natt<br>rustup standard nattlig</p>    Н�n�[ۦ�`�R��b�9ߥ���:�j   
<ol start="0">
<li>./init.sh</li>
<li>skapa api/.env</li>
<li>api/init.sh</li>
<li>api/dev.sh</li>
</ol>
