       )Q���VmV;u�����ͽ8B�	
L| �z   
    O"WeF�DOYp�<����:xz��b��#�Z   <h1>felsökning</h1>
<h2>Installera lokala paket globalt</h2>
<p><code>npm link</code></p>    ��3աb�l��s���:*1vd!)��~�fNWT   
<p>Detta är praktiskt för att felsöka körbara filer i package.json &gt; bin</p>