       ��IJWd��{x�er\���p�)`�ꛯ��  <h2>Försäljningsargument</h2>
<ol start="0">
<li>Fleranvändarbyte utan att logga ut</li>
<li>Internationalisering 121 språk stöds</li>
<li>Separering av främre och bakre ändar</li>
<li>webbkomponent fungerar med alla ramverk</li>
<li>Komponenter kan kombineras efter behag och oanvända främre komponenter stödjer optimering av trädskakning</li>
<li>Stöd för privat driftsättning</li>
<li>Den egenutvecklade verifieringskodmodulen kan även användas i intranätet</li>
<li>Inaktivera engångsregistrering via e-post som standard</li>
<li>Plug-in system, lätt för sekundär utveckling</li>
</ol>
<h2>handledning</h2>
<ol start="0">
<li>Konfigurera användaravtal</li>
</ol>
