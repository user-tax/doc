       )Q���VmV;u�����ͽ8B�	
L| �z   
    8
&)p��4`���|��ݯ�)s���@?��+   <p>last installera sd fd</p>