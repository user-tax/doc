       )Q���VmV;u�����ͽ8B�	
L| �z   
    :�p��%ҡ�(�1؜�	) ���g�C؏��	�   <p><a href="https://user.tax"><img src="https://raw.githubusercontent.com/user-tax/user.tax-img/main/f/logo-txt.svg" alt="Användare. Beskatta" /></a></p>    �G��G��4kͨD���A�����+i���   
<p><a href="https://user-tax.zulipchat.com"><img src="https://raw.githubusercontent.com/user-tax/user.tax-img/main/f/Zulip.svg" alt="Zulip" /></a></p>